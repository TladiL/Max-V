cpu_inst : cpu PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
