c_cpu_inst : c_cpu PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
